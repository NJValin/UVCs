class clk_rstn_cfg extends uvm_object;
	
endclass : clk_rstn_cfg
